module gura

pub const (
	version = '0.1.5'
)
