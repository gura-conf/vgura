module main

import math
import vgura

fn main() {
	data := map{
		'pepe': vgura.Any(math.inf(1))
	}
	text := vgura.encode(data)
	println(text)
}
