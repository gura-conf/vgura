module vgura

pub const (
	version = '0.1.2'
)
